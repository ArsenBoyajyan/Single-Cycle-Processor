module memory(

    );
endmodule
